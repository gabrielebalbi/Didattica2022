
package my_package;

//`ifndef LENGTH
//  `define LENGTH 4   
//`endif

   int unsigned LENGTH = 4;
   
//`include "des_if.sv"
`include "Item.sv"

//`include "scoreboard.sv"
`include "driver.sv"
`include "monitor.sv"
`include "gen_item_seq.sv"
//`include "agent.sv"
//`include "env.sv"
`include "base_test.sv"
//`include "test_1011.sv"

//`define LENGTH 4
//   parameter LENGTH=4;
   
   
endpackage // my_package
   
//import my_package::*;
   
